module control_unit(
	output regDst, 
	output branch,
	output memRead,
	output memWrite,
	output [2:0] ALUop,
	output ALUsrc,
	output regWrite
	output jump,
	output byteOperations,
	output move,

	input [5:0] opcode
);

	//add
	
	//sub
	
	//addi
	
	//subi
	
	//and
	
	//or
	
	//andi
	
	//ori
	
	//lw
	
	//sw
	
	//lb
	
	//sb
	
	//slt
	
	//slti
	
	//beq
	
	//bne
	
	//j
	
	//jal 
	
	//jr
	
	//move
 
endmodule

